
`define cntrl_w(a,b) tb_hydra_lux.odata[a*32+:32]=b;
`define cntrl_r(a,b) b=tb_hydra_lux.idata[a*32+:32];

module hydra_lux_cntrl #(parameter HYDRA_OFFS_O=0,parameter HYDRA_OFFS_I=0)
	();
// input

// conn_file: conn2.txt write
// conn_file: conn0.txt read

// tasks_to_generate
// io_frw_i/hydra/hydra2_0/inst/i_hydra_lux 
	bit [18:0] start_addr; // start_addr[]
	bit [18:0] frame_skip; // frame_skip[]
	bit [7:0] nframes_cyc; // frames_cntr/maxval[] 
	bit   nrst; // ../nrst
	bit stop_nframes; // stop_nframes
	bit [7:2] line_cntv; // line_cntr/val[]
	bit [7:0] frame_cntv; // frames_cntr/val[]
// }
// io_frw_i/hydra/hydra2_0/inst/bramin {
	bit finaddr; // finaddr_reg[]/D
	bit [0:0] stopf; //stopf_reg/D
	bit [11:2] addrb;  // addrb[]
	bit [2:0] ncyc;  // ncyc_reg[]/Q 
	bit ien;  // ien_reg 
// }	
// end_of_tasks_to_generate
/* autogenerated tasks */
task cntrl_w28();
	bit [31:0] odata;
	odata[31:24]=line_cntv[9:2];
	odata[23:16]=frame_cntv[7:0];
	odata[11:0]=addrb[13:2];
	odata[14:12]=ncyc[2:0];
	`cntrl_w(IOCTRL_ADDR_W+28,odata);
endtask;task cntrl_r10();
	bit [31:0] idata;
	`cntrl_r(IOCTRL_ADDR_R+10,idata);
	frame_skip[18:0]=idata[18:0];
	nframes_cyc[7:0]=idata[27:20];
endtask;
task cntrl_r11();
	bit [31:0] idata;
	`cntrl_r(IOCTRL_ADDR_R+11,idata);
	start_addr[18:0]=idata[18:0];
endtask;
task cntrl_r12();
	bit [31:0] idata;
	`cntrl_r(IOCTRL_ADDR_R+12,idata);
	finaddr[11:0]=idata[11:0];
endtask;
/* end autogenerated */
	function [1:0] chr(int bidx); 
		int gn=bidx/6;
		int id=2*(bidx%6);
		chr=chr_concat[gn][id+:2];
	endfunction
	function int chsum(int ch);
		chsum=0;
		//int bidx[2]={24*ch,24*ch+23};
		// wytnij odpowiedni fragment
	endfunction
endmodule	

module deser_la_cntrl #(parameter OFFS_I=0, parameter OFFS_O=0);
	// io_frw_i/lux_in/deser_la_0/inst {
	bit nrst; // nrst
	bit clk_inv; // clk_inv
	bit [1:0] sel1s1; // ch_sel/sel1inst/s1_reg[]/D
	bit [1:0] sel1s2; // ch_sel/sel1inst/s2_reg[]/D
	bit [1:0] sel2s1; // ch_sel/sel2inst/s1_reg[]/D
	bit [1:0] sel2s2; // ch_sel/sel2inst/s2_reg[]/D
	bit [1:0] sel3s1; // ch_sel/sel3inst/s1_reg[]/D
	bit [1:0] sel3s2; // ch_sel/sel3inst/s2_reg[]/D
	//}
// io_frw_i/lux_in/deser_la_0/inst/bramin0 {
	bit [11:0] finaddr; // finaddr_reg[]/D
	bit stopf; //stopf_reg/D
	bit [11:0] addrb;  // addrb[]
	bit [2:0] ncyc;  // ncyc_reg[]/Q 
	bit ien;  // ien_reg 
// }		
// io_frw_i/lux_in/deser_la_0/inst/bramin1 {
	bit [11:0] finaddr1; // finaddr_reg[]/D
	bit stopf1; //stopf_reg/D
	bit [11:0] addrb1;  // addrb[]
	bit [2:0] ncyc1;  // ncyc_reg[]/Q 
	bit ien1;  // ien_reg 
// }		
endmodule	